`timescale 1ns / 1ps



module f(input logic A,B,C,D , output logic Y

    );
    eight_one_mux o1(0,0,0,1,0,1,0,0,1,C,A,Y);
    
endmodule
