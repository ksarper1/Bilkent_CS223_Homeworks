`timescale 1ns / 1ps

module five_thirtytwo_decoder(input [4:0] in, output reg [31:0] ou);
always_comb
    case(in)
                
        0: ou = 32'b00000000000000000000000000000001;
        1: ou = 32'b00000000000000000000000000000010;
        2: ou = 32'b00000000000000000000000000000100;
        3: ou = 32'b00000000000000000000000000001000;
        4: ou = 32'b00000000000000000000000000010000;
        5: ou = 32'b00000000000000000000000000100000;
        6: ou = 32'b00000000000000000000000001000000;
        7: ou = 32'b00000000000000000000000010000000;
        8: ou = 32'b00000000000000000000000100000000;
        9: ou = 32'b00000000000000000000001000000000;
        10: ou = 32'b00000000000000000000010000000000;
        11: ou = 32'b00000000000000000000100000000000;
        12: ou = 32'b00000000000000000001000000000000;
        13: ou = 32'b00000000000000000010000000000000;
        14: ou = 32'b00000000000000000100000000000000;
        15: ou = 32'b00000000000000001000000000000000;
        16: ou = 32'b00000000000000010000000000000000;
        17: ou = 32'b00000000000000100000000000000000;
        18: ou = 32'b00000000000001000000000000000000;
        19: ou = 32'b00000000000010000000000000000000;
        20: ou = 32'b00000000000100000000000000000000;
        21: ou = 32'b00000000001000000000000000000000;
        22: ou = 32'b00000000010000000000000000000000;
        23: ou = 32'b00000000100000000000000000000000;
        24: ou = 32'b00000001000000000000000000000000;
        25: ou = 32'b00000010000000000000000000000000;
        26: ou = 32'b00000100000000000000000000000000;
        27: ou = 32'b00001000000000000000000000000000;
        28: ou = 32'b00010000000000000000000000000000;
        29: ou = 32'b00100000000000000000000000000000;
        30: ou = 32'b01000000000000000000000000000000;
        31: ou = 32'b10000000000000000000000000000000;
        
        
    endcase
endmodule