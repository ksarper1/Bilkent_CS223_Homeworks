`timescale 1ns / 1ps


module four_sixteen_decoder(input [3:0] in, output reg [15:0] ou);
always_comb
    case(in)
                
        0: ou = 16'b0000000000000001;
        1: ou = 16'b0000000000000010;
        2: ou = 16'b0000000000000100;
        3: ou = 16'b0000000000001000;
        4: ou = 16'b0000000000010000;
        5: ou = 16'b0000000000100000;
        6: ou = 16'b0000000001000000;
        7: ou = 16'b0000000010000000;
        8: ou = 16'b0000000100000000;
        9: ou = 16'b0000001000000000;
        10: ou = 16'b0000010000000000;
        11: ou = 16'b0000100000000000;
        12: ou = 16'b0001000000000000;
        13: ou = 16'b0010000000000000;
        14: ou = 16'b0100000000000000;
        15: ou = 16'b1000000000000000;
    endcase
endmodule